`ifndef IP_CONFIG_PKG_SV
 `define IP_CONFIG_PKG_SV

package ip_config_pkg;

   import uvm_pkg::*;      // import the UVM library   
 `include "uvm_macros.svh" // Include the UVM macros

`include "ip_config.sv"


endpackage : ip_config_pkg

`endif